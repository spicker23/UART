module uart();

endmodule
